module problem_7(a, b, c, F);
/* your code below */

endmodule